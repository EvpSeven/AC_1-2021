library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Mux4N is
	generic(N: positive := 32);
	port(in1 	: in std_logic_vector(N-1 downto 0);
		  in2 	: in std_logic_vector(N-1 downto 0);
		  in3 	: in std_logic_vector(N-1 downto 0);
		  in4 	: in std_logic_vector(N-1 downto 0);
		  sel 	: in std_logic_vector(1 downto 0);
		  output : out std_logic_vector(N-1 downto 0));
end MUX4N;

architecture Behavioral of MUX4N is
begin
	process(sel, in1, in2,in3,in4)
	begin
		if(sel = "00") then
			output <= in1;
		elsif( sel = "01") then
			output <= in2;
		elsif(sel = "10") then
			output <= in3;
		elsif(sel = "11") then
			output <= in4;
		end if;
	end process;
end Behavioral;